// nios2_bemicro_system.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module nios2_bemicro_system (
		input  wire        adc_pll_areset_conduit_export,   //   adc_pll_areset_conduit.export
		input  wire [3:0]  button_pio_external_export,      //      button_pio_external.export
		input  wire        clk_clk,                         //                      clk.clk
		inout  wire        i2c_temp_sense_scl_pad_io,       //           i2c_temp_sense.scl_pad_io
		inout  wire        i2c_temp_sense_sda_pad_io,       //                         .sda_pad_io
		output wire [7:0]  led_pio_external_export,         //         led_pio_external.export
		input  wire        reset_reset_n,                   //                    reset.reset_n
		output wire [11:0] sdram_addr,                      //                    sdram.addr
		output wire [1:0]  sdram_ba,                        //                         .ba
		output wire        sdram_cas_n,                     //                         .cas_n
		output wire        sdram_cke,                       //                         .cke
		output wire        sdram_cs_n,                      //                         .cs_n
		inout  wire [15:0] sdram_dq,                        //                         .dq
		output wire [1:0]  sdram_dqm,                       //                         .dqm
		output wire        sdram_ras_n,                     //                         .ras_n
		output wire        sdram_we_n,                      //                         .we_n
		output wire        sdram_pll_80shift_clk,           //        sdram_pll_80shift.clk
		input  wire        sdram_pll_areset_conduit_export, // sdram_pll_areset_conduit.export
		output wire        sdram_pll_locked_conduit_export, // sdram_pll_locked_conduit.export
		input  wire        spi_accelerometer_MISO,          //        spi_accelerometer.MISO
		output wire        spi_accelerometer_MOSI,          //                         .MOSI
		output wire        spi_accelerometer_SCLK,          //                         .SCLK
		output wire        spi_accelerometer_SS_n,          //                         .SS_n
		input  wire        spi_dac_MISO,                    //                  spi_dac.MISO
		output wire        spi_dac_MOSI,                    //                         .MOSI
		output wire        spi_dac_SCLK,                    //                         .SCLK
		output wire        spi_dac_SS_n                     //                         .SS_n
	);

	wire         adc_pll_c0_clk;                                                  // adc_pll:c0 -> modular_adc:adc_pll_clock_clk
	wire         sdram_pll_c0_clk;                                                // sdram_pll:c0 -> [irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, irq_synchronizer_003:sender_clk, mm_interconnect_0:sdram_pll_c0_clk, modular_adc:clock_clk, nios2_cpu:clk, onchip_ram:clk, rst_controller_002:clk, sdram:clk, slow_periph_bridge:s0_clk, spi_accelerometer:clk, spi_dac:clk, ufm_flash:clock]
	wire         sdram_pll_c2_clk;                                                // sdram_pll:c2 -> [button_pio:clk, i2c_temp_sense:wb_clk_i, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, irq_synchronizer_002:receiver_clk, irq_synchronizer_003:receiver_clk, jtag_uart:clk, led_pio:clk, mm_interconnect_1:sdram_pll_c2_clk, rst_controller_001:clk, slow_periph_bridge:m0_clk, sysid:clock, timer:clk]
	wire         adc_pll_locked_conduit_export;                                   // adc_pll:locked -> modular_adc:adc_pll_locked_export
	wire  [31:0] nios2_cpu_data_master_readdata;                                  // mm_interconnect_0:nios2_cpu_data_master_readdata -> nios2_cpu:d_readdata
	wire         nios2_cpu_data_master_waitrequest;                               // mm_interconnect_0:nios2_cpu_data_master_waitrequest -> nios2_cpu:d_waitrequest
	wire         nios2_cpu_data_master_debugaccess;                               // nios2_cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_cpu_data_master_debugaccess
	wire  [25:0] nios2_cpu_data_master_address;                                   // nios2_cpu:d_address -> mm_interconnect_0:nios2_cpu_data_master_address
	wire   [3:0] nios2_cpu_data_master_byteenable;                                // nios2_cpu:d_byteenable -> mm_interconnect_0:nios2_cpu_data_master_byteenable
	wire         nios2_cpu_data_master_read;                                      // nios2_cpu:d_read -> mm_interconnect_0:nios2_cpu_data_master_read
	wire         nios2_cpu_data_master_write;                                     // nios2_cpu:d_write -> mm_interconnect_0:nios2_cpu_data_master_write
	wire  [31:0] nios2_cpu_data_master_writedata;                                 // nios2_cpu:d_writedata -> mm_interconnect_0:nios2_cpu_data_master_writedata
	wire  [31:0] nios2_cpu_instruction_master_readdata;                           // mm_interconnect_0:nios2_cpu_instruction_master_readdata -> nios2_cpu:i_readdata
	wire         nios2_cpu_instruction_master_waitrequest;                        // mm_interconnect_0:nios2_cpu_instruction_master_waitrequest -> nios2_cpu:i_waitrequest
	wire  [25:0] nios2_cpu_instruction_master_address;                            // nios2_cpu:i_address -> mm_interconnect_0:nios2_cpu_instruction_master_address
	wire         nios2_cpu_instruction_master_read;                               // nios2_cpu:i_read -> mm_interconnect_0:nios2_cpu_instruction_master_read
	wire  [31:0] mm_interconnect_0_ufm_flash_csr_readdata;                        // ufm_flash:avmm_csr_readdata -> mm_interconnect_0:ufm_flash_csr_readdata
	wire   [0:0] mm_interconnect_0_ufm_flash_csr_address;                         // mm_interconnect_0:ufm_flash_csr_address -> ufm_flash:avmm_csr_addr
	wire         mm_interconnect_0_ufm_flash_csr_read;                            // mm_interconnect_0:ufm_flash_csr_read -> ufm_flash:avmm_csr_read
	wire         mm_interconnect_0_ufm_flash_csr_write;                           // mm_interconnect_0:ufm_flash_csr_write -> ufm_flash:avmm_csr_write
	wire  [31:0] mm_interconnect_0_ufm_flash_csr_writedata;                       // mm_interconnect_0:ufm_flash_csr_writedata -> ufm_flash:avmm_csr_writedata
	wire  [31:0] mm_interconnect_0_ufm_flash_data_readdata;                       // ufm_flash:avmm_data_readdata -> mm_interconnect_0:ufm_flash_data_readdata
	wire         mm_interconnect_0_ufm_flash_data_waitrequest;                    // ufm_flash:avmm_data_waitrequest -> mm_interconnect_0:ufm_flash_data_waitrequest
	wire  [14:0] mm_interconnect_0_ufm_flash_data_address;                        // mm_interconnect_0:ufm_flash_data_address -> ufm_flash:avmm_data_addr
	wire         mm_interconnect_0_ufm_flash_data_read;                           // mm_interconnect_0:ufm_flash_data_read -> ufm_flash:avmm_data_read
	wire         mm_interconnect_0_ufm_flash_data_readdatavalid;                  // ufm_flash:avmm_data_readdatavalid -> mm_interconnect_0:ufm_flash_data_readdatavalid
	wire         mm_interconnect_0_ufm_flash_data_write;                          // mm_interconnect_0:ufm_flash_data_write -> ufm_flash:avmm_data_write
	wire  [31:0] mm_interconnect_0_ufm_flash_data_writedata;                      // mm_interconnect_0:ufm_flash_data_writedata -> ufm_flash:avmm_data_writedata
	wire   [3:0] mm_interconnect_0_ufm_flash_data_burstcount;                     // mm_interconnect_0:ufm_flash_data_burstcount -> ufm_flash:avmm_data_burstcount
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata;            // nios2_cpu:debug_mem_slave_readdata -> mm_interconnect_0:nios2_cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest;         // nios2_cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:nios2_cpu_debug_mem_slave_debugaccess -> nios2_cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_address;             // mm_interconnect_0:nios2_cpu_debug_mem_slave_address -> nios2_cpu:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_read;                // mm_interconnect_0:nios2_cpu_debug_mem_slave_read -> nios2_cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:nios2_cpu_debug_mem_slave_byteenable -> nios2_cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_write;               // mm_interconnect_0:nios2_cpu_debug_mem_slave_write -> nios2_cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:nios2_cpu_debug_mem_slave_writedata -> nios2_cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_readdata;                  // sdram_pll:readdata -> mm_interconnect_0:sdram_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_sdram_pll_pll_slave_address;                   // mm_interconnect_0:sdram_pll_pll_slave_address -> sdram_pll:address
	wire         mm_interconnect_0_sdram_pll_pll_slave_read;                      // mm_interconnect_0:sdram_pll_pll_slave_read -> sdram_pll:read
	wire         mm_interconnect_0_sdram_pll_pll_slave_write;                     // mm_interconnect_0:sdram_pll_pll_slave_write -> sdram_pll:write
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_writedata;                 // mm_interconnect_0:sdram_pll_pll_slave_writedata -> sdram_pll:writedata
	wire  [31:0] mm_interconnect_0_adc_pll_pll_slave_readdata;                    // adc_pll:readdata -> mm_interconnect_0:adc_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_adc_pll_pll_slave_address;                     // mm_interconnect_0:adc_pll_pll_slave_address -> adc_pll:address
	wire         mm_interconnect_0_adc_pll_pll_slave_read;                        // mm_interconnect_0:adc_pll_pll_slave_read -> adc_pll:read
	wire         mm_interconnect_0_adc_pll_pll_slave_write;                       // mm_interconnect_0:adc_pll_pll_slave_write -> adc_pll:write
	wire  [31:0] mm_interconnect_0_adc_pll_pll_slave_writedata;                   // mm_interconnect_0:adc_pll_pll_slave_writedata -> adc_pll:writedata
	wire  [31:0] mm_interconnect_0_slow_periph_bridge_s0_readdata;                // slow_periph_bridge:s0_readdata -> mm_interconnect_0:slow_periph_bridge_s0_readdata
	wire         mm_interconnect_0_slow_periph_bridge_s0_waitrequest;             // slow_periph_bridge:s0_waitrequest -> mm_interconnect_0:slow_periph_bridge_s0_waitrequest
	wire         mm_interconnect_0_slow_periph_bridge_s0_debugaccess;             // mm_interconnect_0:slow_periph_bridge_s0_debugaccess -> slow_periph_bridge:s0_debugaccess
	wire   [9:0] mm_interconnect_0_slow_periph_bridge_s0_address;                 // mm_interconnect_0:slow_periph_bridge_s0_address -> slow_periph_bridge:s0_address
	wire         mm_interconnect_0_slow_periph_bridge_s0_read;                    // mm_interconnect_0:slow_periph_bridge_s0_read -> slow_periph_bridge:s0_read
	wire   [3:0] mm_interconnect_0_slow_periph_bridge_s0_byteenable;              // mm_interconnect_0:slow_periph_bridge_s0_byteenable -> slow_periph_bridge:s0_byteenable
	wire         mm_interconnect_0_slow_periph_bridge_s0_readdatavalid;           // slow_periph_bridge:s0_readdatavalid -> mm_interconnect_0:slow_periph_bridge_s0_readdatavalid
	wire         mm_interconnect_0_slow_periph_bridge_s0_write;                   // mm_interconnect_0:slow_periph_bridge_s0_write -> slow_periph_bridge:s0_write
	wire  [31:0] mm_interconnect_0_slow_periph_bridge_s0_writedata;               // mm_interconnect_0:slow_periph_bridge_s0_writedata -> slow_periph_bridge:s0_writedata
	wire   [0:0] mm_interconnect_0_slow_periph_bridge_s0_burstcount;              // mm_interconnect_0:slow_periph_bridge_s0_burstcount -> slow_periph_bridge:s0_burstcount
	wire         mm_interconnect_0_onchip_ram_s1_chipselect;                      // mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_readdata;                        // onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_ram_s1_address;                         // mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	wire   [3:0] mm_interconnect_0_onchip_ram_s1_byteenable;                      // mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	wire         mm_interconnect_0_onchip_ram_s1_write;                           // mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_writedata;                       // mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	wire         mm_interconnect_0_onchip_ram_s1_clken;                           // mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                           // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                             // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                          // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [21:0] mm_interconnect_0_sdram_s1_address;                              // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                 // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                           // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                        // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                            // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [31:0] mm_interconnect_0_modular_adc_sample_store_csr_readdata;         // modular_adc:sample_store_csr_readdata -> mm_interconnect_0:modular_adc_sample_store_csr_readdata
	wire   [6:0] mm_interconnect_0_modular_adc_sample_store_csr_address;          // mm_interconnect_0:modular_adc_sample_store_csr_address -> modular_adc:sample_store_csr_address
	wire         mm_interconnect_0_modular_adc_sample_store_csr_read;             // mm_interconnect_0:modular_adc_sample_store_csr_read -> modular_adc:sample_store_csr_read
	wire         mm_interconnect_0_modular_adc_sample_store_csr_write;            // mm_interconnect_0:modular_adc_sample_store_csr_write -> modular_adc:sample_store_csr_write
	wire  [31:0] mm_interconnect_0_modular_adc_sample_store_csr_writedata;        // mm_interconnect_0:modular_adc_sample_store_csr_writedata -> modular_adc:sample_store_csr_writedata
	wire  [31:0] mm_interconnect_0_modular_adc_sequencer_csr_readdata;            // modular_adc:sequencer_csr_readdata -> mm_interconnect_0:modular_adc_sequencer_csr_readdata
	wire   [0:0] mm_interconnect_0_modular_adc_sequencer_csr_address;             // mm_interconnect_0:modular_adc_sequencer_csr_address -> modular_adc:sequencer_csr_address
	wire         mm_interconnect_0_modular_adc_sequencer_csr_read;                // mm_interconnect_0:modular_adc_sequencer_csr_read -> modular_adc:sequencer_csr_read
	wire         mm_interconnect_0_modular_adc_sequencer_csr_write;               // mm_interconnect_0:modular_adc_sequencer_csr_write -> modular_adc:sequencer_csr_write
	wire  [31:0] mm_interconnect_0_modular_adc_sequencer_csr_writedata;           // mm_interconnect_0:modular_adc_sequencer_csr_writedata -> modular_adc:sequencer_csr_writedata
	wire         mm_interconnect_0_spi_accelerometer_spi_control_port_chipselect; // mm_interconnect_0:spi_accelerometer_spi_control_port_chipselect -> spi_accelerometer:spi_select
	wire  [15:0] mm_interconnect_0_spi_accelerometer_spi_control_port_readdata;   // spi_accelerometer:data_to_cpu -> mm_interconnect_0:spi_accelerometer_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_accelerometer_spi_control_port_address;    // mm_interconnect_0:spi_accelerometer_spi_control_port_address -> spi_accelerometer:mem_addr
	wire         mm_interconnect_0_spi_accelerometer_spi_control_port_read;       // mm_interconnect_0:spi_accelerometer_spi_control_port_read -> spi_accelerometer:read_n
	wire         mm_interconnect_0_spi_accelerometer_spi_control_port_write;      // mm_interconnect_0:spi_accelerometer_spi_control_port_write -> spi_accelerometer:write_n
	wire  [15:0] mm_interconnect_0_spi_accelerometer_spi_control_port_writedata;  // mm_interconnect_0:spi_accelerometer_spi_control_port_writedata -> spi_accelerometer:data_from_cpu
	wire         mm_interconnect_0_spi_dac_spi_control_port_chipselect;           // mm_interconnect_0:spi_dac_spi_control_port_chipselect -> spi_dac:spi_select
	wire  [15:0] mm_interconnect_0_spi_dac_spi_control_port_readdata;             // spi_dac:data_to_cpu -> mm_interconnect_0:spi_dac_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_dac_spi_control_port_address;              // mm_interconnect_0:spi_dac_spi_control_port_address -> spi_dac:mem_addr
	wire         mm_interconnect_0_spi_dac_spi_control_port_read;                 // mm_interconnect_0:spi_dac_spi_control_port_read -> spi_dac:read_n
	wire         mm_interconnect_0_spi_dac_spi_control_port_write;                // mm_interconnect_0:spi_dac_spi_control_port_write -> spi_dac:write_n
	wire  [15:0] mm_interconnect_0_spi_dac_spi_control_port_writedata;            // mm_interconnect_0:spi_dac_spi_control_port_writedata -> spi_dac:data_from_cpu
	wire         slow_periph_bridge_m0_waitrequest;                               // mm_interconnect_1:slow_periph_bridge_m0_waitrequest -> slow_periph_bridge:m0_waitrequest
	wire  [31:0] slow_periph_bridge_m0_readdata;                                  // mm_interconnect_1:slow_periph_bridge_m0_readdata -> slow_periph_bridge:m0_readdata
	wire         slow_periph_bridge_m0_debugaccess;                               // slow_periph_bridge:m0_debugaccess -> mm_interconnect_1:slow_periph_bridge_m0_debugaccess
	wire   [9:0] slow_periph_bridge_m0_address;                                   // slow_periph_bridge:m0_address -> mm_interconnect_1:slow_periph_bridge_m0_address
	wire         slow_periph_bridge_m0_read;                                      // slow_periph_bridge:m0_read -> mm_interconnect_1:slow_periph_bridge_m0_read
	wire   [3:0] slow_periph_bridge_m0_byteenable;                                // slow_periph_bridge:m0_byteenable -> mm_interconnect_1:slow_periph_bridge_m0_byteenable
	wire         slow_periph_bridge_m0_readdatavalid;                             // mm_interconnect_1:slow_periph_bridge_m0_readdatavalid -> slow_periph_bridge:m0_readdatavalid
	wire  [31:0] slow_periph_bridge_m0_writedata;                                 // slow_periph_bridge:m0_writedata -> mm_interconnect_1:slow_periph_bridge_m0_writedata
	wire         slow_periph_bridge_m0_write;                                     // slow_periph_bridge:m0_write -> mm_interconnect_1:slow_periph_bridge_m0_write
	wire   [0:0] slow_periph_bridge_m0_burstcount;                                // slow_periph_bridge:m0_burstcount -> mm_interconnect_1:slow_periph_bridge_m0_burstcount
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;        // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;          // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest;       // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;           // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;              // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;             // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;         // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_1_i2c_temp_sense_avalon_slave_0_chipselect;      // mm_interconnect_1:i2c_temp_sense_avalon_slave_0_chipselect -> i2c_temp_sense:wb_stb_i
	wire   [7:0] mm_interconnect_1_i2c_temp_sense_avalon_slave_0_readdata;        // i2c_temp_sense:wb_dat_o -> mm_interconnect_1:i2c_temp_sense_avalon_slave_0_readdata
	wire         mm_interconnect_1_i2c_temp_sense_avalon_slave_0_waitrequest;     // i2c_temp_sense:wb_ack_o -> mm_interconnect_1:i2c_temp_sense_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_1_i2c_temp_sense_avalon_slave_0_address;         // mm_interconnect_1:i2c_temp_sense_avalon_slave_0_address -> i2c_temp_sense:wb_adr_i
	wire         mm_interconnect_1_i2c_temp_sense_avalon_slave_0_write;           // mm_interconnect_1:i2c_temp_sense_avalon_slave_0_write -> i2c_temp_sense:wb_we_i
	wire   [7:0] mm_interconnect_1_i2c_temp_sense_avalon_slave_0_writedata;       // mm_interconnect_1:i2c_temp_sense_avalon_slave_0_writedata -> i2c_temp_sense:wb_dat_i
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;                  // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;                   // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire         mm_interconnect_1_led_pio_s1_chipselect;                         // mm_interconnect_1:led_pio_s1_chipselect -> led_pio:chipselect
	wire  [31:0] mm_interconnect_1_led_pio_s1_readdata;                           // led_pio:readdata -> mm_interconnect_1:led_pio_s1_readdata
	wire   [1:0] mm_interconnect_1_led_pio_s1_address;                            // mm_interconnect_1:led_pio_s1_address -> led_pio:address
	wire         mm_interconnect_1_led_pio_s1_write;                              // mm_interconnect_1:led_pio_s1_write -> led_pio:write_n
	wire  [31:0] mm_interconnect_1_led_pio_s1_writedata;                          // mm_interconnect_1:led_pio_s1_writedata -> led_pio:writedata
	wire         mm_interconnect_1_button_pio_s1_chipselect;                      // mm_interconnect_1:button_pio_s1_chipselect -> button_pio:chipselect
	wire  [31:0] mm_interconnect_1_button_pio_s1_readdata;                        // button_pio:readdata -> mm_interconnect_1:button_pio_s1_readdata
	wire   [1:0] mm_interconnect_1_button_pio_s1_address;                         // mm_interconnect_1:button_pio_s1_address -> button_pio:address
	wire         mm_interconnect_1_button_pio_s1_write;                           // mm_interconnect_1:button_pio_s1_write -> button_pio:write_n
	wire  [31:0] mm_interconnect_1_button_pio_s1_writedata;                       // mm_interconnect_1:button_pio_s1_writedata -> button_pio:writedata
	wire         mm_interconnect_1_timer_s1_chipselect;                           // mm_interconnect_1:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_1_timer_s1_readdata;                             // timer:readdata -> mm_interconnect_1:timer_s1_readdata
	wire   [2:0] mm_interconnect_1_timer_s1_address;                              // mm_interconnect_1:timer_s1_address -> timer:address
	wire         mm_interconnect_1_timer_s1_write;                                // mm_interconnect_1:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_1_timer_s1_writedata;                            // mm_interconnect_1:timer_s1_writedata -> timer:writedata
	wire         irq_mapper_receiver1_irq;                                        // spi_accelerometer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                        // spi_dac:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver6_irq;                                        // modular_adc:sample_store_irq_irq -> irq_mapper:receiver6_irq
	wire  [31:0] nios2_cpu_irq_irq;                                               // irq_mapper:sender_irq -> nios2_cpu:irq
	wire         irq_mapper_receiver0_irq;                                        // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                   // i2c_temp_sense:wb_inta_o -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver3_irq;                                        // irq_synchronizer_001:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                               // jtag_uart:av_irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver4_irq;                                        // irq_synchronizer_002:sender_irq -> irq_mapper:receiver4_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                               // timer:irq -> irq_synchronizer_002:receiver_irq
	wire         irq_mapper_receiver5_irq;                                        // irq_synchronizer_003:sender_irq -> irq_mapper:receiver5_irq
	wire   [0:0] irq_synchronizer_003_receiver_irq;                               // button_pio:irq -> irq_synchronizer_003:receiver_irq
	wire         rst_controller_reset_out_reset;                                  // rst_controller:reset_out -> [adc_pll:reset, mm_interconnect_0:sdram_pll_inclk_interface_reset_reset_bridge_in_reset_reset, sdram_pll:reset]
	wire         nios2_cpu_debug_reset_request_reset;                             // nios2_cpu:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;                              // rst_controller_001:reset_out -> [button_pio:reset_n, i2c_temp_sense:wb_rst_i, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, jtag_uart:rst_n, led_pio:reset_n, mm_interconnect_1:slow_periph_bridge_m0_reset_reset_bridge_in_reset_reset, slow_periph_bridge:m0_reset, sysid:reset_n, timer:reset_n]
	wire         rst_controller_002_reset_out_reset;                              // rst_controller_002:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, mm_interconnect_0:nios2_cpu_reset_reset_bridge_in_reset_reset, modular_adc:reset_sink_reset_n, nios2_cpu:reset_n, onchip_ram:reset, rst_translator:in_reset, sdram:reset_n, slow_periph_bridge:s0_reset, spi_accelerometer:reset_n, spi_dac:reset_n, ufm_flash:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                          // rst_controller_002:reset_req -> [nios2_cpu:reset_req, onchip_ram:reset_req, rst_translator:reset_req_in]

	nios2_bemicro_system_adc_pll adc_pll (
		.clk                (clk_clk),                                       //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                // inclk_interface_reset.reset
		.read               (mm_interconnect_0_adc_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_adc_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_adc_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_adc_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_adc_pll_pll_slave_writedata), //                      .writedata
		.c0                 (adc_pll_c0_clk),                                //                    c0.clk
		.areset             (adc_pll_areset_conduit_export),                 //        areset_conduit.export
		.locked             (adc_pll_locked_conduit_export),                 //        locked_conduit.export
		.phasedone          (),                                              //           (terminated)
		.phasecounterselect (3'b000),                                        //           (terminated)
		.phaseupdown        (1'b0),                                          //           (terminated)
		.phasestep          (1'b0),                                          //           (terminated)
		.scanclk            (1'b0)                                           //           (terminated)
	);

	nios2_bemicro_system_button_pio button_pio (
		.clk        (sdram_pll_c2_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_1_button_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_button_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_button_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_button_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_button_pio_s1_readdata),   //                    .readdata
		.in_port    (button_pio_external_export),                 // external_connection.export
		.irq        (irq_synchronizer_003_receiver_irq)           //                 irq.irq
	);

	i2c_opencores i2c_temp_sense (
		.wb_clk_i   (sdram_pll_c2_clk),                                            //            clock.clk
		.wb_rst_i   (rst_controller_001_reset_out_reset),                          //      clock_reset.reset
		.scl_pad_io (i2c_temp_sense_scl_pad_io),                                   //           export.export
		.sda_pad_io (i2c_temp_sense_sda_pad_io),                                   //                 .export
		.wb_adr_i   (mm_interconnect_1_i2c_temp_sense_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_1_i2c_temp_sense_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_1_i2c_temp_sense_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_1_i2c_temp_sense_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_1_i2c_temp_sense_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_1_i2c_temp_sense_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_synchronizer_receiver_irq)                                // interrupt_sender.irq
	);

	nios2_bemicro_system_jtag_uart jtag_uart (
		.clk            (sdram_pll_c2_clk),                                          //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_001_receiver_irq)                          //               irq.irq
	);

	nios2_bemicro_system_led_pio led_pio (
		.clk        (sdram_pll_c2_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_pio_s1_readdata),   //                    .readdata
		.out_port   (led_pio_external_export)                  // external_connection.export
	);

	nios2_bemicro_system_modular_adc modular_adc (
		.clock_clk                  (sdram_pll_c0_clk),                                         //            clock.clk
		.reset_sink_reset_n         (~rst_controller_002_reset_out_reset),                      //       reset_sink.reset_n
		.adc_pll_clock_clk          (adc_pll_c0_clk),                                           //    adc_pll_clock.clk
		.adc_pll_locked_export      (adc_pll_locked_conduit_export),                            //   adc_pll_locked.export
		.sequencer_csr_address      (mm_interconnect_0_modular_adc_sequencer_csr_address),      //    sequencer_csr.address
		.sequencer_csr_read         (mm_interconnect_0_modular_adc_sequencer_csr_read),         //                 .read
		.sequencer_csr_write        (mm_interconnect_0_modular_adc_sequencer_csr_write),        //                 .write
		.sequencer_csr_writedata    (mm_interconnect_0_modular_adc_sequencer_csr_writedata),    //                 .writedata
		.sequencer_csr_readdata     (mm_interconnect_0_modular_adc_sequencer_csr_readdata),     //                 .readdata
		.sample_store_csr_address   (mm_interconnect_0_modular_adc_sample_store_csr_address),   // sample_store_csr.address
		.sample_store_csr_read      (mm_interconnect_0_modular_adc_sample_store_csr_read),      //                 .read
		.sample_store_csr_write     (mm_interconnect_0_modular_adc_sample_store_csr_write),     //                 .write
		.sample_store_csr_writedata (mm_interconnect_0_modular_adc_sample_store_csr_writedata), //                 .writedata
		.sample_store_csr_readdata  (mm_interconnect_0_modular_adc_sample_store_csr_readdata),  //                 .readdata
		.sample_store_irq_irq       (irq_mapper_receiver6_irq)                                  // sample_store_irq.irq
	);

	nios2_bemicro_system_nios2_cpu nios2_cpu (
		.clk                                 (sdram_pll_c0_clk),                                        //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_cpu_data_master_read),                              //                          .read
		.d_readdata                          (nios2_cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_cpu_data_master_write),                             //                          .write
		.d_writedata                         (nios2_cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                         // custom_instruction_master.readra
	);

	nios2_bemicro_system_onchip_ram onchip_ram (
		.clk        (sdram_pll_c0_clk),                           //   clk1.clk
		.address    (mm_interconnect_0_onchip_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req)      //       .reset_req
	);

	nios2_bemicro_system_sdram sdram (
		.clk            (sdram_pll_c0_clk),                         //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	nios2_bemicro_system_sdram_pll sdram_pll (
		.clk                (clk_clk),                                         //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                  // inclk_interface_reset.reset
		.read               (mm_interconnect_0_sdram_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_sdram_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_sdram_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_sdram_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_sdram_pll_pll_slave_writedata), //                      .writedata
		.c0                 (sdram_pll_c0_clk),                                //                    c0.clk
		.c1                 (sdram_pll_80shift_clk),                           //                    c1.clk
		.c2                 (sdram_pll_c2_clk),                                //                    c2.clk
		.areset             (sdram_pll_areset_conduit_export),                 //        areset_conduit.export
		.locked             (sdram_pll_locked_conduit_export),                 //        locked_conduit.export
		.phasedone          (),                                                //           (terminated)
		.phasecounterselect (3'b000),                                          //           (terminated)
		.phaseupdown        (1'b0),                                            //           (terminated)
		.phasestep          (1'b0),                                            //           (terminated)
		.scanclk            (1'b0)                                             //           (terminated)
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (32),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) slow_periph_bridge (
		.m0_clk           (sdram_pll_c2_clk),                                      //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                    // m0_reset.reset
		.s0_clk           (sdram_pll_c0_clk),                                      //   s0_clk.clk
		.s0_reset         (rst_controller_002_reset_out_reset),                    // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_slow_periph_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_slow_periph_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_slow_periph_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_slow_periph_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_slow_periph_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_slow_periph_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_slow_periph_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_slow_periph_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_slow_periph_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_slow_periph_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (slow_periph_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (slow_periph_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (slow_periph_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (slow_periph_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (slow_periph_bridge_m0_writedata),                       //         .writedata
		.m0_address       (slow_periph_bridge_m0_address),                         //         .address
		.m0_write         (slow_periph_bridge_m0_write),                           //         .write
		.m0_read          (slow_periph_bridge_m0_read),                            //         .read
		.m0_byteenable    (slow_periph_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (slow_periph_bridge_m0_debugaccess)                      //         .debugaccess
	);

	nios2_bemicro_system_spi_accelerometer spi_accelerometer (
		.clk           (sdram_pll_c0_clk),                                                //              clk.clk
		.reset_n       (~rst_controller_002_reset_out_reset),                             //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_accelerometer_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_accelerometer_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_accelerometer_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_accelerometer_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_accelerometer_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_accelerometer_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver1_irq),                                        //              irq.irq
		.MISO          (spi_accelerometer_MISO),                                          //         external.export
		.MOSI          (spi_accelerometer_MOSI),                                          //                 .export
		.SCLK          (spi_accelerometer_SCLK),                                          //                 .export
		.SS_n          (spi_accelerometer_SS_n)                                           //                 .export
	);

	nios2_bemicro_system_spi_accelerometer spi_dac (
		.clk           (sdram_pll_c0_clk),                                      //              clk.clk
		.reset_n       (~rst_controller_002_reset_out_reset),                   //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_dac_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_dac_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_dac_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_dac_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_dac_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_dac_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver2_irq),                              //              irq.irq
		.MISO          (spi_dac_MISO),                                          //         external.export
		.MOSI          (spi_dac_MOSI),                                          //                 .export
		.SCLK          (spi_dac_SCLK),                                          //                 .export
		.SS_n          (spi_dac_SS_n)                                           //                 .export
	);

	nios2_bemicro_system_sysid sysid (
		.clock    (sdram_pll_c2_clk),                               //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	nios2_bemicro_system_timer timer (
		.clk        (sdram_pll_c2_clk),                      //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_1_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_002_receiver_irq)      //   irq.irq
	);

	altera_onchip_flash #(
		.INIT_FILENAME                       (""),
		.INIT_FILENAME_SIM                   (""),
		.DEVICE_FAMILY                       ("MAX 10"),
		.PART_NAME                           ("10M08DAF484C8GES"),
		.DEVICE_ID                           ("08"),
		.SECTOR1_START_ADDR                  (0),
		.SECTOR1_END_ADDR                    (4095),
		.SECTOR2_START_ADDR                  (4096),
		.SECTOR2_END_ADDR                    (8191),
		.SECTOR3_START_ADDR                  (8192),
		.SECTOR3_END_ADDR                    (29183),
		.SECTOR4_START_ADDR                  (0),
		.SECTOR4_END_ADDR                    (0),
		.SECTOR5_START_ADDR                  (0),
		.SECTOR5_END_ADDR                    (0),
		.MIN_VALID_ADDR                      (0),
		.MAX_VALID_ADDR                      (29183),
		.MIN_UFM_VALID_ADDR                  (0),
		.MAX_UFM_VALID_ADDR                  (29183),
		.SECTOR1_MAP                         (1),
		.SECTOR2_MAP                         (2),
		.SECTOR3_MAP                         (3),
		.SECTOR4_MAP                         (0),
		.SECTOR5_MAP                         (0),
		.ADDR_RANGE1_END_ADDR                (29183),
		.ADDR_RANGE1_OFFSET                  (512),
		.ADDR_RANGE2_OFFSET                  (0),
		.AVMM_DATA_ADDR_WIDTH                (15),
		.AVMM_DATA_DATA_WIDTH                (32),
		.AVMM_DATA_BURSTCOUNT_WIDTH          (4),
		.SECTOR_READ_PROTECTION_MODE         (28),
		.FLASH_SEQ_READ_DATA_COUNT           (2),
		.FLASH_ADDR_ALIGNMENT_BITS           (1),
		.FLASH_READ_CYCLE_MAX_INDEX          (4),
		.FLASH_RESET_CYCLE_MAX_INDEX         (20),
		.FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  (96),
		.FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX (28000000),
		.FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX (24400),
		.PARALLEL_MODE                       (1),
		.READ_AND_WRITE_MODE                 (1),
		.WRAPPING_BURST_MODE                 (0),
		.IS_DUAL_BOOT                        ("False"),
		.IS_ERAM_SKIP                        ("True"),
		.IS_COMPRESSED_IMAGE                 ("False")
	) ufm_flash (
		.clock                   (sdram_pll_c0_clk),                               //    clk.clk
		.reset_n                 (~rst_controller_002_reset_out_reset),            // nreset.reset_n
		.avmm_data_addr          (mm_interconnect_0_ufm_flash_data_address),       //   data.address
		.avmm_data_read          (mm_interconnect_0_ufm_flash_data_read),          //       .read
		.avmm_data_writedata     (mm_interconnect_0_ufm_flash_data_writedata),     //       .writedata
		.avmm_data_write         (mm_interconnect_0_ufm_flash_data_write),         //       .write
		.avmm_data_readdata      (mm_interconnect_0_ufm_flash_data_readdata),      //       .readdata
		.avmm_data_waitrequest   (mm_interconnect_0_ufm_flash_data_waitrequest),   //       .waitrequest
		.avmm_data_readdatavalid (mm_interconnect_0_ufm_flash_data_readdatavalid), //       .readdatavalid
		.avmm_data_burstcount    (mm_interconnect_0_ufm_flash_data_burstcount),    //       .burstcount
		.avmm_csr_addr           (mm_interconnect_0_ufm_flash_csr_address),        //    csr.address
		.avmm_csr_read           (mm_interconnect_0_ufm_flash_csr_read),           //       .read
		.avmm_csr_writedata      (mm_interconnect_0_ufm_flash_csr_writedata),      //       .writedata
		.avmm_csr_write          (mm_interconnect_0_ufm_flash_csr_write),          //       .write
		.avmm_csr_readdata       (mm_interconnect_0_ufm_flash_csr_readdata)        //       .readdata
	);

	nios2_bemicro_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                               (clk_clk),                                                         //                                             clk_0_clk.clk
		.sdram_pll_c0_clk                                            (sdram_pll_c0_clk),                                                //                                          sdram_pll_c0.clk
		.nios2_cpu_reset_reset_bridge_in_reset_reset                 (rst_controller_002_reset_out_reset),                              //                 nios2_cpu_reset_reset_bridge_in_reset.reset
		.sdram_pll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                  // sdram_pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.nios2_cpu_data_master_address                               (nios2_cpu_data_master_address),                                   //                                 nios2_cpu_data_master.address
		.nios2_cpu_data_master_waitrequest                           (nios2_cpu_data_master_waitrequest),                               //                                                      .waitrequest
		.nios2_cpu_data_master_byteenable                            (nios2_cpu_data_master_byteenable),                                //                                                      .byteenable
		.nios2_cpu_data_master_read                                  (nios2_cpu_data_master_read),                                      //                                                      .read
		.nios2_cpu_data_master_readdata                              (nios2_cpu_data_master_readdata),                                  //                                                      .readdata
		.nios2_cpu_data_master_write                                 (nios2_cpu_data_master_write),                                     //                                                      .write
		.nios2_cpu_data_master_writedata                             (nios2_cpu_data_master_writedata),                                 //                                                      .writedata
		.nios2_cpu_data_master_debugaccess                           (nios2_cpu_data_master_debugaccess),                               //                                                      .debugaccess
		.nios2_cpu_instruction_master_address                        (nios2_cpu_instruction_master_address),                            //                          nios2_cpu_instruction_master.address
		.nios2_cpu_instruction_master_waitrequest                    (nios2_cpu_instruction_master_waitrequest),                        //                                                      .waitrequest
		.nios2_cpu_instruction_master_read                           (nios2_cpu_instruction_master_read),                               //                                                      .read
		.nios2_cpu_instruction_master_readdata                       (nios2_cpu_instruction_master_readdata),                           //                                                      .readdata
		.adc_pll_pll_slave_address                                   (mm_interconnect_0_adc_pll_pll_slave_address),                     //                                     adc_pll_pll_slave.address
		.adc_pll_pll_slave_write                                     (mm_interconnect_0_adc_pll_pll_slave_write),                       //                                                      .write
		.adc_pll_pll_slave_read                                      (mm_interconnect_0_adc_pll_pll_slave_read),                        //                                                      .read
		.adc_pll_pll_slave_readdata                                  (mm_interconnect_0_adc_pll_pll_slave_readdata),                    //                                                      .readdata
		.adc_pll_pll_slave_writedata                                 (mm_interconnect_0_adc_pll_pll_slave_writedata),                   //                                                      .writedata
		.modular_adc_sample_store_csr_address                        (mm_interconnect_0_modular_adc_sample_store_csr_address),          //                          modular_adc_sample_store_csr.address
		.modular_adc_sample_store_csr_write                          (mm_interconnect_0_modular_adc_sample_store_csr_write),            //                                                      .write
		.modular_adc_sample_store_csr_read                           (mm_interconnect_0_modular_adc_sample_store_csr_read),             //                                                      .read
		.modular_adc_sample_store_csr_readdata                       (mm_interconnect_0_modular_adc_sample_store_csr_readdata),         //                                                      .readdata
		.modular_adc_sample_store_csr_writedata                      (mm_interconnect_0_modular_adc_sample_store_csr_writedata),        //                                                      .writedata
		.modular_adc_sequencer_csr_address                           (mm_interconnect_0_modular_adc_sequencer_csr_address),             //                             modular_adc_sequencer_csr.address
		.modular_adc_sequencer_csr_write                             (mm_interconnect_0_modular_adc_sequencer_csr_write),               //                                                      .write
		.modular_adc_sequencer_csr_read                              (mm_interconnect_0_modular_adc_sequencer_csr_read),                //                                                      .read
		.modular_adc_sequencer_csr_readdata                          (mm_interconnect_0_modular_adc_sequencer_csr_readdata),            //                                                      .readdata
		.modular_adc_sequencer_csr_writedata                         (mm_interconnect_0_modular_adc_sequencer_csr_writedata),           //                                                      .writedata
		.nios2_cpu_debug_mem_slave_address                           (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),             //                             nios2_cpu_debug_mem_slave.address
		.nios2_cpu_debug_mem_slave_write                             (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),               //                                                      .write
		.nios2_cpu_debug_mem_slave_read                              (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),                //                                                      .read
		.nios2_cpu_debug_mem_slave_readdata                          (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),            //                                                      .readdata
		.nios2_cpu_debug_mem_slave_writedata                         (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),           //                                                      .writedata
		.nios2_cpu_debug_mem_slave_byteenable                        (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),          //                                                      .byteenable
		.nios2_cpu_debug_mem_slave_waitrequest                       (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest),         //                                                      .waitrequest
		.nios2_cpu_debug_mem_slave_debugaccess                       (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess),         //                                                      .debugaccess
		.onchip_ram_s1_address                                       (mm_interconnect_0_onchip_ram_s1_address),                         //                                         onchip_ram_s1.address
		.onchip_ram_s1_write                                         (mm_interconnect_0_onchip_ram_s1_write),                           //                                                      .write
		.onchip_ram_s1_readdata                                      (mm_interconnect_0_onchip_ram_s1_readdata),                        //                                                      .readdata
		.onchip_ram_s1_writedata                                     (mm_interconnect_0_onchip_ram_s1_writedata),                       //                                                      .writedata
		.onchip_ram_s1_byteenable                                    (mm_interconnect_0_onchip_ram_s1_byteenable),                      //                                                      .byteenable
		.onchip_ram_s1_chipselect                                    (mm_interconnect_0_onchip_ram_s1_chipselect),                      //                                                      .chipselect
		.onchip_ram_s1_clken                                         (mm_interconnect_0_onchip_ram_s1_clken),                           //                                                      .clken
		.sdram_s1_address                                            (mm_interconnect_0_sdram_s1_address),                              //                                              sdram_s1.address
		.sdram_s1_write                                              (mm_interconnect_0_sdram_s1_write),                                //                                                      .write
		.sdram_s1_read                                               (mm_interconnect_0_sdram_s1_read),                                 //                                                      .read
		.sdram_s1_readdata                                           (mm_interconnect_0_sdram_s1_readdata),                             //                                                      .readdata
		.sdram_s1_writedata                                          (mm_interconnect_0_sdram_s1_writedata),                            //                                                      .writedata
		.sdram_s1_byteenable                                         (mm_interconnect_0_sdram_s1_byteenable),                           //                                                      .byteenable
		.sdram_s1_readdatavalid                                      (mm_interconnect_0_sdram_s1_readdatavalid),                        //                                                      .readdatavalid
		.sdram_s1_waitrequest                                        (mm_interconnect_0_sdram_s1_waitrequest),                          //                                                      .waitrequest
		.sdram_s1_chipselect                                         (mm_interconnect_0_sdram_s1_chipselect),                           //                                                      .chipselect
		.sdram_pll_pll_slave_address                                 (mm_interconnect_0_sdram_pll_pll_slave_address),                   //                                   sdram_pll_pll_slave.address
		.sdram_pll_pll_slave_write                                   (mm_interconnect_0_sdram_pll_pll_slave_write),                     //                                                      .write
		.sdram_pll_pll_slave_read                                    (mm_interconnect_0_sdram_pll_pll_slave_read),                      //                                                      .read
		.sdram_pll_pll_slave_readdata                                (mm_interconnect_0_sdram_pll_pll_slave_readdata),                  //                                                      .readdata
		.sdram_pll_pll_slave_writedata                               (mm_interconnect_0_sdram_pll_pll_slave_writedata),                 //                                                      .writedata
		.slow_periph_bridge_s0_address                               (mm_interconnect_0_slow_periph_bridge_s0_address),                 //                                 slow_periph_bridge_s0.address
		.slow_periph_bridge_s0_write                                 (mm_interconnect_0_slow_periph_bridge_s0_write),                   //                                                      .write
		.slow_periph_bridge_s0_read                                  (mm_interconnect_0_slow_periph_bridge_s0_read),                    //                                                      .read
		.slow_periph_bridge_s0_readdata                              (mm_interconnect_0_slow_periph_bridge_s0_readdata),                //                                                      .readdata
		.slow_periph_bridge_s0_writedata                             (mm_interconnect_0_slow_periph_bridge_s0_writedata),               //                                                      .writedata
		.slow_periph_bridge_s0_burstcount                            (mm_interconnect_0_slow_periph_bridge_s0_burstcount),              //                                                      .burstcount
		.slow_periph_bridge_s0_byteenable                            (mm_interconnect_0_slow_periph_bridge_s0_byteenable),              //                                                      .byteenable
		.slow_periph_bridge_s0_readdatavalid                         (mm_interconnect_0_slow_periph_bridge_s0_readdatavalid),           //                                                      .readdatavalid
		.slow_periph_bridge_s0_waitrequest                           (mm_interconnect_0_slow_periph_bridge_s0_waitrequest),             //                                                      .waitrequest
		.slow_periph_bridge_s0_debugaccess                           (mm_interconnect_0_slow_periph_bridge_s0_debugaccess),             //                                                      .debugaccess
		.spi_accelerometer_spi_control_port_address                  (mm_interconnect_0_spi_accelerometer_spi_control_port_address),    //                    spi_accelerometer_spi_control_port.address
		.spi_accelerometer_spi_control_port_write                    (mm_interconnect_0_spi_accelerometer_spi_control_port_write),      //                                                      .write
		.spi_accelerometer_spi_control_port_read                     (mm_interconnect_0_spi_accelerometer_spi_control_port_read),       //                                                      .read
		.spi_accelerometer_spi_control_port_readdata                 (mm_interconnect_0_spi_accelerometer_spi_control_port_readdata),   //                                                      .readdata
		.spi_accelerometer_spi_control_port_writedata                (mm_interconnect_0_spi_accelerometer_spi_control_port_writedata),  //                                                      .writedata
		.spi_accelerometer_spi_control_port_chipselect               (mm_interconnect_0_spi_accelerometer_spi_control_port_chipselect), //                                                      .chipselect
		.spi_dac_spi_control_port_address                            (mm_interconnect_0_spi_dac_spi_control_port_address),              //                              spi_dac_spi_control_port.address
		.spi_dac_spi_control_port_write                              (mm_interconnect_0_spi_dac_spi_control_port_write),                //                                                      .write
		.spi_dac_spi_control_port_read                               (mm_interconnect_0_spi_dac_spi_control_port_read),                 //                                                      .read
		.spi_dac_spi_control_port_readdata                           (mm_interconnect_0_spi_dac_spi_control_port_readdata),             //                                                      .readdata
		.spi_dac_spi_control_port_writedata                          (mm_interconnect_0_spi_dac_spi_control_port_writedata),            //                                                      .writedata
		.spi_dac_spi_control_port_chipselect                         (mm_interconnect_0_spi_dac_spi_control_port_chipselect),           //                                                      .chipselect
		.ufm_flash_csr_address                                       (mm_interconnect_0_ufm_flash_csr_address),                         //                                         ufm_flash_csr.address
		.ufm_flash_csr_write                                         (mm_interconnect_0_ufm_flash_csr_write),                           //                                                      .write
		.ufm_flash_csr_read                                          (mm_interconnect_0_ufm_flash_csr_read),                            //                                                      .read
		.ufm_flash_csr_readdata                                      (mm_interconnect_0_ufm_flash_csr_readdata),                        //                                                      .readdata
		.ufm_flash_csr_writedata                                     (mm_interconnect_0_ufm_flash_csr_writedata),                       //                                                      .writedata
		.ufm_flash_data_address                                      (mm_interconnect_0_ufm_flash_data_address),                        //                                        ufm_flash_data.address
		.ufm_flash_data_write                                        (mm_interconnect_0_ufm_flash_data_write),                          //                                                      .write
		.ufm_flash_data_read                                         (mm_interconnect_0_ufm_flash_data_read),                           //                                                      .read
		.ufm_flash_data_readdata                                     (mm_interconnect_0_ufm_flash_data_readdata),                       //                                                      .readdata
		.ufm_flash_data_writedata                                    (mm_interconnect_0_ufm_flash_data_writedata),                      //                                                      .writedata
		.ufm_flash_data_burstcount                                   (mm_interconnect_0_ufm_flash_data_burstcount),                     //                                                      .burstcount
		.ufm_flash_data_readdatavalid                                (mm_interconnect_0_ufm_flash_data_readdatavalid),                  //                                                      .readdatavalid
		.ufm_flash_data_waitrequest                                  (mm_interconnect_0_ufm_flash_data_waitrequest)                     //                                                      .waitrequest
	);

	nios2_bemicro_system_mm_interconnect_1 mm_interconnect_1 (
		.sdram_pll_c2_clk                                        (sdram_pll_c2_clk),                                             //                                      sdram_pll_c2.clk
		.slow_periph_bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                           // slow_periph_bridge_m0_reset_reset_bridge_in_reset.reset
		.slow_periph_bridge_m0_address                           (slow_periph_bridge_m0_address),                                //                             slow_periph_bridge_m0.address
		.slow_periph_bridge_m0_waitrequest                       (slow_periph_bridge_m0_waitrequest),                            //                                                  .waitrequest
		.slow_periph_bridge_m0_burstcount                        (slow_periph_bridge_m0_burstcount),                             //                                                  .burstcount
		.slow_periph_bridge_m0_byteenable                        (slow_periph_bridge_m0_byteenable),                             //                                                  .byteenable
		.slow_periph_bridge_m0_read                              (slow_periph_bridge_m0_read),                                   //                                                  .read
		.slow_periph_bridge_m0_readdata                          (slow_periph_bridge_m0_readdata),                               //                                                  .readdata
		.slow_periph_bridge_m0_readdatavalid                     (slow_periph_bridge_m0_readdatavalid),                          //                                                  .readdatavalid
		.slow_periph_bridge_m0_write                             (slow_periph_bridge_m0_write),                                  //                                                  .write
		.slow_periph_bridge_m0_writedata                         (slow_periph_bridge_m0_writedata),                              //                                                  .writedata
		.slow_periph_bridge_m0_debugaccess                       (slow_periph_bridge_m0_debugaccess),                            //                                                  .debugaccess
		.button_pio_s1_address                                   (mm_interconnect_1_button_pio_s1_address),                      //                                     button_pio_s1.address
		.button_pio_s1_write                                     (mm_interconnect_1_button_pio_s1_write),                        //                                                  .write
		.button_pio_s1_readdata                                  (mm_interconnect_1_button_pio_s1_readdata),                     //                                                  .readdata
		.button_pio_s1_writedata                                 (mm_interconnect_1_button_pio_s1_writedata),                    //                                                  .writedata
		.button_pio_s1_chipselect                                (mm_interconnect_1_button_pio_s1_chipselect),                   //                                                  .chipselect
		.i2c_temp_sense_avalon_slave_0_address                   (mm_interconnect_1_i2c_temp_sense_avalon_slave_0_address),      //                     i2c_temp_sense_avalon_slave_0.address
		.i2c_temp_sense_avalon_slave_0_write                     (mm_interconnect_1_i2c_temp_sense_avalon_slave_0_write),        //                                                  .write
		.i2c_temp_sense_avalon_slave_0_readdata                  (mm_interconnect_1_i2c_temp_sense_avalon_slave_0_readdata),     //                                                  .readdata
		.i2c_temp_sense_avalon_slave_0_writedata                 (mm_interconnect_1_i2c_temp_sense_avalon_slave_0_writedata),    //                                                  .writedata
		.i2c_temp_sense_avalon_slave_0_waitrequest               (~mm_interconnect_1_i2c_temp_sense_avalon_slave_0_waitrequest), //                                                  .waitrequest
		.i2c_temp_sense_avalon_slave_0_chipselect                (mm_interconnect_1_i2c_temp_sense_avalon_slave_0_chipselect),   //                                                  .chipselect
		.jtag_uart_avalon_jtag_slave_address                     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),        //                       jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                       (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),          //                                                  .write
		.jtag_uart_avalon_jtag_slave_read                        (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),           //                                                  .read
		.jtag_uart_avalon_jtag_slave_readdata                    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),       //                                                  .readdata
		.jtag_uart_avalon_jtag_slave_writedata                   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),      //                                                  .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                 (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest),    //                                                  .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),     //                                                  .chipselect
		.led_pio_s1_address                                      (mm_interconnect_1_led_pio_s1_address),                         //                                        led_pio_s1.address
		.led_pio_s1_write                                        (mm_interconnect_1_led_pio_s1_write),                           //                                                  .write
		.led_pio_s1_readdata                                     (mm_interconnect_1_led_pio_s1_readdata),                        //                                                  .readdata
		.led_pio_s1_writedata                                    (mm_interconnect_1_led_pio_s1_writedata),                       //                                                  .writedata
		.led_pio_s1_chipselect                                   (mm_interconnect_1_led_pio_s1_chipselect),                      //                                                  .chipselect
		.sysid_control_slave_address                             (mm_interconnect_1_sysid_control_slave_address),                //                               sysid_control_slave.address
		.sysid_control_slave_readdata                            (mm_interconnect_1_sysid_control_slave_readdata),               //                                                  .readdata
		.timer_s1_address                                        (mm_interconnect_1_timer_s1_address),                           //                                          timer_s1.address
		.timer_s1_write                                          (mm_interconnect_1_timer_s1_write),                             //                                                  .write
		.timer_s1_readdata                                       (mm_interconnect_1_timer_s1_readdata),                          //                                                  .readdata
		.timer_s1_writedata                                      (mm_interconnect_1_timer_s1_writedata),                         //                                                  .writedata
		.timer_s1_chipselect                                     (mm_interconnect_1_timer_s1_chipselect)                         //                                                  .chipselect
	);

	nios2_bemicro_system_irq_mapper irq_mapper (
		.clk           (sdram_pll_c0_clk),                   //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),           // receiver6.irq
		.sender_irq    (nios2_cpu_irq_irq)                   //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (sdram_pll_c2_clk),                   //       receiver_clk.clk
		.sender_clk     (sdram_pll_c0_clk),                   //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (sdram_pll_c2_clk),                   //       receiver_clk.clk
		.sender_clk     (sdram_pll_c0_clk),                   //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (sdram_pll_c2_clk),                   //       receiver_clk.clk
		.sender_clk     (sdram_pll_c0_clk),                   //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (sdram_pll_c2_clk),                   //       receiver_clk.clk
		.sender_clk     (sdram_pll_c0_clk),                   //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver5_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (nios2_cpu_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (nios2_cpu_debug_reset_request_reset), // reset_in1.reset
		.clk            (sdram_pll_c2_clk),                    //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_cpu_debug_reset_request_reset),    // reset_in1.reset
		.clk            (sdram_pll_c0_clk),                       //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
